r65c02_rom_32768words_8bits_inst : r65c02_rom_32768words_8bits PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		rden	 => rden_sig,
		q	 => q_sig
	);
